(** This module implements a signature *)
Module Type Signature.

Parameter Kappa:Type.
Parameter Arity:Kappa-> nat.

End Signature.

Print Signature.